library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


entity clk_digital is
	port(
		clk_40 			: in std_logic;
		hpos    			: in integer;
		vpos				: in integer;
		videoOn			: in std_logic;
		GPIO_0         : in std_logic_vector(3 downto 0);
		clk_low        : in std_logic;
	   cntr59         : in integer;
		cntr59_min     : in integer;
		cntr59_hour    : in integer;
		
		--outputs
		VGA_R          : out std_logic_vector(9 downto 0);
		VGA_G          : out std_logic_vector(9 downto 0);
		VGA_B          : out std_logic_vector(9 downto 0)
	);
end entity;


architecture clk_digital of clk_digital is

	signal cntr59_hour_sig : integer;
		
	signal vpos1_dig: integer:=0;
	signal hpos1_dig: integer:=0;
	signal vpos2_dig: integer:=0;
	signal hpos2_dig: integer:=0;
	

	signal ycoord_init_dig: integer:=320;
	signal ycoord_end_dig : integer:=400;
	signal xcoord_init_dig: integer:=200;
	signal xcoord_end_dig : integer:=600;
	
	
	signal VGA_R_sig : std_logic_vector(9 downto 0);
	signal VGA_G_sig : std_logic_vector(9 downto 0);
	signal VGA_B_sig : std_logic_vector(9 downto 0);
		
	type HFZ_dig is array (0 to 79) of std_logic_vector(0 to 39);
								
constant BM_0_dig: HFZ_dig :=("0000000000000000000000000000000000000000",--1
								      "0000000000000000000000000000000000000000",--2
								      "0011111111111111111111111111111111111100",--3
								      "0011111111111111111111111111111111111100",--4
									   "0011111111111111111111111111111111111100",--5
									   "0011111111111111111111111111111111111100",--6
									   "0011111111111111111111111111111111111100",--7
									   "0011111111111111111111111111111111111100",--8
									   "0011111111111111111111111111111111111100",--9
								      "0011111111111111111111111111111111111100",--10         --0
								      "0011111111000000000000000000001111111100",--11
								      "0011111111000000000000000000001111111100",--12
								      "0011111111000000000000000000001111111100",--13
								      "0011111111000000000000000000001111111100",--14
								      "0011111111000000000000000000001111111100",--15
								      "0011111111000000000000000000001111111100",--16
								      "0011111111000000000000000000001111111100",--17
								      "0011111111000000000000000000001111111100",--18
								      "0011111111000000000000000000001111111100",--19
								      "0011111111000000000000000000001111111100",     --20
									   "0011111111000000000000000000001111111100",--1
								      "0011111111000000000000000000001111111100",--2
								      "0011111111000000000000000000001111111100",--3
								      "0011111111000000000000000000001111111100",--4
									   "0011111111000000000000000000001111111100",--5
									   "0011111111000000000000000000001111111100",--6
									   "0011111111000000000000000000001111111100",--7
									   "0011111111000000000000000000001111111100",--8
									   "0011111111000000000000000000001111111100",--9
								      "0011111111000000000000000000001111111100",--10         --0
								      "0011111111000000000000000000001111111100",--11
								      "0011111111000000000000000000001111111100",--12
								      "0011111111000000000000000000001111111100",--13
								      "0011111111000000000000000000001111111100",--14
								      "0011111111000000000000000000001111111100",--15
								      "0011111111000000000000000000001111111100",--16
								      "0011111111000000000000000000001111111100",--17
								      "0011111111000000000000000000001111111100",--18
								      "0011111111000000000000000000001111111100",--19
								      "0011111111000000000000000000001111111100",     --40
									   "0011111111000000000000000000001111111100",--1
								      "0011111111000000000000000000001111111100",--2
								      "0011111111000000000000000000001111111100",--3
								      "0011111111000000000000000000001111111100",--4
									   "0011111111000000000000000000001111111100",--5
									   "0011111111000000000000000000001111111100",--6
									   "0011111111000000000000000000001111111100",--7
									   "0011111111000000000000000000001111111100",--8
									   "0011111111000000000000000000001111111100",--9
								      "0011111111000000000000000000001111111100",--10         --0
								      "0011111111000000000000000000001111111100",--11
								      "0011111111000000000000000000001111111100",--12
								      "0011111111000000000000000000001111111100",--13
								      "0011111111000000000000000000001111111100",--14
								      "0011111111000000000000000000001111111100",--15
								      "0011111111000000000000000000001111111100",--16
								      "0011111111000000000000000000001111111100",--17
								      "0011111111000000000000000000001111111100",--18
								      "0011111111000000000000000000001111111100",--19
								      "0011111111000000000000000000001111111100",    --60
									   "0011111111000000000000000000001111111100",--1
								      "0011111111000000000000000000001111111100",--2
								      "0011111111000000000000000000001111111100",--3
								      "0011111111000000000000000000001111111100",--4
									   "0011111111000000000000000000001111111100",--5
									   "0011111111000000000000000000001111111100",--6
									   "0011111111000000000000000000001111111100",--7
									   "0011111111000000000000000000001111111100",--8
									   "0011111111000000000000000000001111111100",--9
								      "0011111111000000000000000000001111111100",--10         --0
								      "0011111111111111111111111111111111111100",--11
								      "0011111111111111111111111111111111111100",--12
								      "0011111111111111111111111111111111111100",--13
								      "0011111111111111111111111111111111111100",--14
								      "0011111111111111111111111111111111111100",--15
								      "0011111111111111111111111111111111111100",--16
								      "0011111111111111111111111111111111111100",--17
								      "0011111111111111111111111111111111111100",--18
								      "0000000000000000000000000000000000000000",--19
								      "0000000000000000000000000000000000000000");  --80
									 
	   constant BM_BOS_dig:HFZ_dig:=("0000000000000000000000000000000000000000",--1
								            "0000000000000000000000000000000000000000",--2
								            "0000000000000000000000000000000000000000",--3  
								            "0000000000000000000000000000000000000000",--4
									         "0000000000000000000000000000000000000000",--5
									         "0000000000000000000000000000000000000000",--6
									         "0000000000000000000000000000000000000000",--7
									         "0000000000000000000000000000000000000000",--8
									         "0000000000000000000000000000000000000000",--9
								            "0000000000000000000000000000000000000000",--10         --BOS
								            "0000000000000000000000000000000000000000",--11
								            "0000000000000000000000000000000000000000",--12
								            "0000000000000000000000000000000000000000",--13
								            "0000000000000000000000000000000000000000",--14
								            "0000000000000000000000000000000000000000",--15
								            "0000000000000000000000000000000000000000",--16
								            "0000000000000000000000000000000000000000",--17
								            "0000000000000000000000000000000000000000",--18
								            "0000000000000000000000000000000000000000",--19
								            "0000000000000000000000000000000000000000",     --20
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000",
									         "0000000000000000000000000000000000000000");
									 
										 
									 
									 
	   constant BM_1_dig:HFZ_dig:=  ("0000000000000000000000000000000000000000",--1
								    "0000000000000000000000000000000011111110",--2
								    "0000000000000000000000000000000011111110",--3
								    "0000000000000000000000000000000011111110",--4
									 "0000000000000000000000000000000011111110",--5
									 "0000000000000000000000000000000011111110",--6
									 "0000000000000000000000000000000011111110",--7
									 "0000000000000000000000000000000011111110",--8
									 "0000000000000000000000000000000011111110",--9
								    "0000000000000000000000000000000011111110",--10         --1
								    "0000000000000000000000000000000011111110",--11
								    "0000000000000000000000000000000011111110",--12
								    "0000000000000000000000000000000011111110",--13
								    "0000000000000000000000000000000011111110",--14
								    "0000000000000000000000000000000011111110",--15
								    "0000000000000000000000000000000011111110",--16
								    "0000000000000000000000000000000011111110",--17
								    "0000000000000000000000000000000011111110",--18
								    "0000000000000000000000000000000011111110",--19
								    "0000000000000000000000000000000011111110",     --20
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000011111110",
									 "0000000000000000000000000000000000000000");	
									 
	  constant BM_2_dig: HFZ_dig :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0111111111111111111111111111111111111110",--6
									 "0111111111111111111111111111111111111110",--7
									 "0111111111111111111111111111111111111110",--8
									 "0111111111111111111111111111111111111110",--9
								    "0000000000000000000000000000000111111110",--10         --22222222222
								    "0000000000000000000000000000000111111110",--11                  --222222222222
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0000000000000000000000000000000111111110",--17
								    "0000000000000000000000000000000111111110",--18
								    "0000000000000000000000000000000111111110",--19
								    "0000000000000000000000000000000111111110",     --20
									 "0000000000000000000000000000000111111110",--1
								    "0000000000000000000000000000000111111110",--2
								    "0000000000000000000000000000000111111110",--3
								    "0000000000000000000000000000000111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111110000000000000000000000000000000",--5
									 "0111111110000000000000000000000000000000",--6
									 "0111111110000000000000000000000000000000",--7
									 "0111111110000000000000000000000000000000",--8
									 "0111111110000000000000000000000000000000",--9
								    "0111111110000000000000000000000000000000",--10         
								    "0111111110000000000000000000000000000000",--11
								    "0111111110000000000000000000000000000000",--12
								    "0111111110000000000000000000000000000000",--13
								    "0111111110000000000000000000000000000000",--14
								    "0111111110000000000000000000000000000000",--15
								    "0111111110000000000000000000000000000000",--16
								    "0111111110000000000000000000000000000000",--17
								    "0111111110000000000000000000000000000000",--18
								    "0111111110000000000000000000000000000000",--19
								    "0111111110000000000000000000000000000000",    --60
									 "0111111110000000000000000000000000000000",--1
								    "0111111110000000000000000000000000000000",--2
								    "0111111110000000000000000000000000000000",--3
								    "0111111110000000000000000000000000000000",--4
									 "0111111110000000000000000000000000000000",--5
									 "0111111110000000000000000000000000000000",--6
									 "0111111110000000000000000000000000000000",--7
									 "0111111110000000000000000000000000000000",--8
									 "0111111110000000000000000000000000000000",--9
								    "0111111110000000000000000000000000000000",--10         
								    "0111111110000000000000000000000000000000",--11
								    "0111111111111111111111111111111111111110",--12
								    "0111111111111111111111111111111111111110",--13
								    "0111111111111111111111111111111111111110",--14
								    "0111111111111111111111111111111111111110",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80

		  constant BM_3_dig: HFZ_dig :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0111111111111111111111111111111111111110",--6
									 "0111111111111111111111111111111111111110",--7
									 "0111111111111111111111111111111111111110",--8
									 "0111111111111111111111111111111111111110",--9
								    "0000000000000000000000000000000111111110",--10         --33333333
								    "0000000000000000000000000000000111111110",--11                
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0000000000000000000000000000000111111110",--17
								    "0000000000000000000000000000000111111110",--18
								    "0000000000000000000000000000000111111110",--19
								    "0000000000000000000000000000000111111110",     --20
									 "0000000000000000000000000000000111111110",--1
								    "0000000000000000000000000000000111111110",--2
								    "0000000000000000000000000000000111111110",--3
								    "0000000000000000000000000000000111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0000000000000000000000000000000111111110",--17
								    "0000000000000000000000000000000111111110",--18
								    "0000000000000000000000000000000111111110",--19
								    "0000000000000000000000000000000111111110",    --60
									 "0000000000000000000000000000000111111110",--1
								    "0000000000000000000000000000000111111110",--2
								    "0000000000000000000000000000000111111110",--3
								    "0000000000000000000000000000000111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0111111111111111111111111111111111111110",--12
								    "0111111111111111111111111111111111111110",--13
								    "0111111111111111111111111111111111111110",--14
								    "0111111111111111111111111111111111111110",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
		
		constant BM_4_dig: HFZ_dig :=("0000000000000000000000000000000000000000",--1
								    "0111111110000000000000000000000111111110",--2
								    "0111111110000000000000000000000111111110",--3
								    "0111111110000000000000000000000111111110",--4
									 "0111111110000000000000000000000111111110",--5
									 "0111111110000000000000000000000111111110",--6
									 "0111111110000000000000000000000111111110",--7
									 "0111111110000000000000000000000111111110",--8
									 "0111111110000000000000000000000111111110",--9
								    "0111111110000000000000000000000111111110",--10         --4
								    "0111111110000000000000000000000111111110",--11                
								    "0111111110000000000000000000000111111110",--12
								    "0111111110000000000000000000000111111110",--13
								    "0111111110000000000000000000000111111110",--14
								    "0111111110000000000000000000000111111110",--15
								    "0111111110000000000000000000000111111110",--16
								    "0111111110000000000000000000000111111110",--17
								    "0111111110000000000000000000000111111110",--18
								    "0111111110000000000000000000000111111110",--19
								    "0111111110000000000000000000000111111110",     --20
									 "0111111110000000000000000000000111111110",--1
								    "0111111110000000000000000000000111111110",--2
								    "0111111110000000000000000000000111111110",--3
								    "0111111110000000000000000000000111111110",--4
									 "0111111110000000000000000000000111111110",--5
									 "0111111110000000000000000000000111111110",--6
									 "0111111110000000000000000000000111111110",--7
									 "0111111110000000000000000000000111111110",--8
									 "0111111110000000000000000000000111111110",--9
								    "0111111110000000000000000000000111111110",--10         
								    "0111111110000000000000000000000111111110",--11
								    "0111111110000000000000000000000111111110",--12
								    "0111111110000000000000000000000111111110",--13
								    "0111111110000000000000000000000111111110",--14
								    "0111111110000000000000000000000111111110",--15
								    "0111111110000000000000000000000111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0000000000000000000000000000000111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0000000000000000000000000000000111111110",--17
								    "0000000000000000000000000000000111111110",--18
								    "0000000000000000000000000000000111111110",--19
								    "0000000000000000000000000000000111111110",    --60
									 "0000000000000000000000000000000111111110",--1
								    "0000000000000000000000000000000111111110",--2
								    "0000000000000000000000000000000111111110",--3
								    "0000000000000000000000000000000111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0000000000000000000000000000000111111110",--17
								    "0000000000000000000000000000000111111110",--18
								    "0000000000000000000000000000000111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
									 
									 
      constant BM_5_dig: HFZ_dig :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0111111111111111111111111111111111111110",--6
									 "0111111111111111111111111111111111111110",--7
									 "0111111111111111111111111111111111111110",--8
									 "0111111111111111111111111111111111111110",--9
								    "0111111110000000000000000000000000000000",--10         
								    "0111111110000000000000000000000000000000",--11                  --5
								    "0111111110000000000000000000000000000000",--12
								    "0111111110000000000000000000000000000000",--13
								    "0111111110000000000000000000000000000000",--14
								    "0111111110000000000000000000000000000000",--15
								    "0111111110000000000000000000000000000000",--16
								    "0111111110000000000000000000000000000000",--17
								    "0111111110000000000000000000000000000000",--18
								    "0111111110000000000000000000000000000000",--19
								    "0111111110000000000000000000000000000000",     --20
									 "0111111110000000000000000000000000000000",--1
								    "0111111110000000000000000000000000000000",--2
								    "0111111110000000000000000000000000000000",--3
								    "0111111110000000000000000000000000000000",--4
									 "0111111110000000000000000000000000000000",--5
									 "0111111110000000000000000000000000000000",--6
									 "0111111110000000000000000000000000000000",--7
									 "0111111110000000000000000000000000000000",--8
									 "0111111110000000000000000000000000000000",--9
								    "0111111110000000000000000000000000000000",--10         
								    "0111111110000000000000000000000000000000",--11
								    "0111111110000000000000000000000000000000",--12
								    "0111111110000000000000000000000000000000",--13
								    "0111111110000000000000000000000000000000",--14
								    "0111111110000000000000000000000000000000",--15
								    "0111111110000000000000000000000000000000",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0000000000000000000000000000000111111110",--17
								    "0000000000000000000000000000000111111110",--18
								    "0000000000000000000000000000000111111110",--19
								    "0000000000000000000000000000000111111110",    --60
									 "0000000000000000000000000000000111111110",--1
								    "0000000000000000000000000000000111111110",--2
								    "0000000000000000000000000000000111111110",--3
								    "0000000000000000000000000000000111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0111111111111111111111111111111111111110",--12
								    "0111111111111111111111111111111111111110",--13
								    "0111111111111111111111111111111111111110",--14
								    "0111111111111111111111111111111111111110",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
									 
      constant BM_6_dig: HFZ_dig :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0111111111111111111111111111111111111110",--6
									 "0111111111111111111111111111111111111110",--7
									 "0111111111111111111111111111111111111100",--8
									 "0111111111111111111111111111111111111100",--9
								    "0111111110000000000000000000000000000000",--10         --6
								    "0111111110000000000000000000000000000000",--11              
								    "0111111110000000000000000000000000000000",--12
								    "0111111110000000000000000000000000000000",--13
								    "0111111110000000000000000000000000000000",--14
								    "0111111110000000000000000000000000000000",--15
								    "0111111110000000000000000000000000000000",--16
								    "0111111110000000000000000000000000000000",--17
								    "0111111110000000000000000000000000000000",--18
								    "0111111110000000000000000000000000000000",--19
								    "0111111110000000000000000000000000000000",     --20
									 "0111111110000000000000000000000000000000",--1
								    "0111111110000000000000000000000000000000",--2
								    "0111111110000000000000000000000000000000",--3
								    "0111111110000000000000000000000000000000",--4
									 "0111111110000000000000000000000000000000",--5
									 "0111111110000000000000000000000000000000",--6
									 "0111111110000000000000000000000000000000",--7
									 "0111111110000000000000000000000000000000",--8
									 "0111111110000000000000000000000000000000",--9
								    "0111111110000000000000000000000000000000",--10         
								    "0111111110000000000000000000000000000000",--11
								    "0111111110000000000000000000000000000000",--12
								    "0111111110000000000000000000000000000000",--13
								    "0111111110000000000000000000000000000000",--14
								    "0111111110000000000000000000000000000000",--15
								    "0111111110000000000000000000000000000000",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111110000000000000000000000111111110",--5
									 "0111111110000000000000000000000111111110",--6
									 "0111111110000000000000000000000111111110",--7
									 "0111111110000000000000000000000111111110",--8
									 "0111111110000000000000000000000111111110",--9
								    "0111111110000000000000000000000111111110",--10         
								    "0111111110000000000000000000000111111110",--11
								    "0111111110000000000000000000000111111110",--12
								    "0111111110000000000000000000000111111110",--13
								    "0111111110000000000000000000000111111110",--14
								    "0111111110000000000000000000000111111110",--15
								    "0111111110000000000000000000000111111110",--16
								    "0111111110000000000000000000000111111110",--17
								    "0111111110000000000000000000000111111110",--18
								    "0111111110000000000000000000000111111110",--19
								    "0111111110000000000000000000000111111110",    --60
									 "0111111110000000000000000000000111111110",--1
								    "0111111110000000000000000000000111111110",--2
								    "0111111110000000000000000000000111111110",--3
								    "0111111110000000000000000000000111111110",--4
									 "0111111110000000000000000000000111111110",--5
									 "0111111110000000000000000000000111111110",--6
									 "0111111110000000000000000000000111111110",--7
									 "0111111110000000000000000000000111111110",--8
									 "0111111110000000000000000000000111111110",--9
								    "0111111110000000000000000000000111111110",--10         
								    "0111111110000000000000000000000111111110",--11
								    "0111111111111111111111111111111111111110",--12
								    "0111111111111111111111111111111111111110",--13
								    "0111111111111111111111111111111111111110",--14
								    "0111111111111111111111111111111111111110",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
									 
	   constant BM_7_dig: HFZ_dig :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0111111111111111111111111111111111111110",--6
									 "0111111111111111111111111111111111111110",--7
									 "0111111111111111111111111111111111111110",--8
									 "0111111111111111111111111111111111111110",--9
								    "0000000000000000000000000000000111111110",--10         --7
								    "0000000000000000000000000000000111111110",--11                
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0000000000000000000000000000000111111110",--17
								    "0000000000000000000000000000000111111110",--18
								    "0000000000000000000000000000000111111110",--19
								    "0000000000000000000000000000000111111110",     --20
									 "0000000000000000000000000000000111111110",--1
								    "0000000000000000000000000000000111111110",--2
								    "0000000000000000000000000000000111111110",--3
								    "0000000000000000000000000000000111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0000000000000000000000000000000111111110",--17
								    "0000000000000000000000000000000111111110",--18
								    "0000000000000000000000000000000111111110",--19
								    "0000000000000000000000000000000111111110",     --40
									 "0000000000000000000000000000000111111110",--1
								    "0000000000000000000000000000000111111110",--2
								    "0000000000000000000000000000000111111110",--3
								    "0000000000000000000000000000000111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0000000000000000000000000000000111111110",--17
								    "0000000000000000000000000000000111111110",--18
								    "0000000000000000000000000000000111111110",--19
								    "0000000000000000000000000000000111111110",    --60
									 "0000000000000000000000000000000111111110",--1
								    "0000000000000000000000000000000111111110",--2
								    "0000000000000000000000000000000111111110",--3
								    "0000000000000000000000000000000111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0000000000000000000000000000000111111110",--17
								    "0000000000000000000000000000000111111110",--18
								    "0000000000000000000000000000000111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
	   constant BM_8_dig: HFZ_dig :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0111111111111111111111111111111111111110",--6
									 "0111111111111111111111111111111111111110",--7
									 "0111111111111111111111111111111111111110",--8
									 "0111111111111111111111111111111111111110",--9
								    "0111111110000000000000000000000111111110",--10         
								    "0111111110000000000000000000000111111110",--11                  --8
								    "0111111110000000000000000000000111111110",--12
								    "0111111110000000000000000000000111111110",--13
								    "0111111110000000000000000000000111111110",--14
								    "0111111110000000000000000000000111111110",--15
								    "0111111110000000000000000000000111111110",--16
								    "0111111110000000000000000000000111111110",--17
								    "0111111110000000000000000000000111111110",--18
								    "0111111110000000000000000000000111111110",--19
								    "0111111110000000000000000000000111111110",     --20
									 "0111111110000000000000000000000111111110",--1
								    "0111111110000000000000000000000111111110",--2
								    "0111111110000000000000000000000111111110",--3
								    "0111111110000000000000000000000111111110",--4
									 "0111111110000000000000000000000111111110",--5
									 "0111111110000000000000000000000111111110",--6
									 "0111111110000000000000000000000111111110",--7
									 "0111111110000000000000000000000111111110",--8
									 "0111111110000000000000000000000111111110",--9
								    "0111111110000000000000000000000111111110",--10         
								    "0111111110000000000000000000000111111110",--11
								    "0111111110000000000000000000000111111110",--12
								    "0111111110000000000000000000000111111110",--13
								    "0111111110000000000000000000000111111110",--14
								    "0111111110000000000000000000000111111110",--15
								    "0111111110000000000000000000000111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111110000000000000000000000111111110",--5
									 "0111111110000000000000000000000111111110",--6
									 "0111111110000000000000000000000111111110",--7
									 "0111111110000000000000000000000111111110",--8
									 "0111111110000000000000000000000111111110",--9
								    "0111111110000000000000000000000111111110",--10         
								    "0111111110000000000000000000000111111110",--11
								    "0111111110000000000000000000000111111110",--12
								    "0111111110000000000000000000000111111110",--13
								    "0111111110000000000000000000000111111110",--14
								    "0111111110000000000000000000000111111110",--15
								    "0111111110000000000000000000000111111110",--16
								    "0111111110000000000000000000000111111110",--17
								    "0111111110000000000000000000000111111110",--18
								    "0111111110000000000000000000000111111110",--19
								    "0111111110000000000000000000000111111110",    --60
									 "0111111110000000000000000000000111111110",--1
								    "0111111110000000000000000000000111111110",--2
								    "0111111110000000000000000000000111111110",--3
								    "0111111110000000000000000000000111111110",--4
									 "0111111110000000000000000000000111111110",--5
									 "0111111110000000000000000000000111111110",--6
									 "0111111110000000000000000000000111111110",--7
									 "0111111110000000000000000000000111111110",--8
									 "0111111110000000000000000000000111111110",--9
								    "0111111110000000000000000000000111111110",--10         
								    "0111111110000000000000000000000111111110",--11
								    "0111111111111111111111111111111111111110",--12
								    "0111111111111111111111111111111111111110",--13
								    "0111111111111111111111111111111111111110",--14
								    "0111111111111111111111111111111111111110",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
									 
	   constant BM_9_dig: HFZ_dig :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0111111111111111111111111111111111111110",--6
									 "0111111111111111111111111111111111111110",--7
									 "0111111111111111111111111111111111111110",--8
									 "0111111111111111111111111111111111111110",--9
								    "0111111110000000000000000000000111111110",--10         
								    "0111111110000000000000000000000111111110",--11                  --9
								    "0111111110000000000000000000000111111110",--12
								    "0111111110000000000000000000000111111110",--13
								    "0111111110000000000000000000000111111110",--14
								    "0111111110000000000000000000000111111110",--15
								    "0111111110000000000000000000000111111110",--16
								    "0111111110000000000000000000000111111110",--17
								    "0111111110000000000000000000000111111110",--18
								    "0111111110000000000000000000000111111110",--19
								    "0111111110000000000000000000000111111110",     --20
									 "0111111110000000000000000000000111111110",--1
								    "0111111110000000000000000000000111111110",--2
								    "0111111110000000000000000000000111111110",--3
								    "0111111110000000000000000000000111111110",--4
									 "0111111110000000000000000000000111111110",--5
									 "0111111110000000000000000000000111111110",--6
									 "0111111110000000000000000000000111111110",--7
									 "0111111110000000000000000000000111111110",--8
									 "0111111110000000000000000000000111111110",--9
								    "0111111110000000000000000000000111111110",--10         
								    "0111111110000000000000000000000111111110",--11
								    "0111111110000000000000000000000111111110",--12
								    "0111111110000000000000000000000111111110",--13
								    "0111111110000000000000000000000111111110",--14
								    "0111111110000000000000000000000111111110",--15
								    "0111111110000000000000000000000111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0000000000000000000000000000000111111110",--12
								    "0000000000000000000000000000000111111110",--13
								    "0000000000000000000000000000000111111110",--14
								    "0000000000000000000000000000000111111110",--15
								    "0000000000000000000000000000000111111110",--16
								    "0000000000000000000000000000000111111110",--17
								    "0000000000000000000000000000000111111110",--18
								    "0000000000000000000000000000000111111110",--19
								    "0000000000000000000000000000000111111110",    --60
									 "0000000000000000000000000000000111111110",--1
								    "0000000000000000000000000000000111111110",--2
								    "0000000000000000000000000000000111111110",--3
								    "0000000000000000000000000000000111111110",--4
									 "0000000000000000000000000000000111111110",--5
									 "0000000000000000000000000000000111111110",--6
									 "0000000000000000000000000000000111111110",--7
									 "0000000000000000000000000000000111111110",--8
									 "0000000000000000000000000000000111111110",--9
								    "0000000000000000000000000000000111111110",--10         
								    "0000000000000000000000000000000111111110",--11
								    "0111111111111111111111111111111111111110",--12
								    "0111111111111111111111111111111111111110",--13
								    "0111111111111111111111111111111111111110",--14
								    "0111111111111111111111111111111111111110",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 

								

									 
	
constant BM_iki_nokta_dig:HFZ_dig:=("0000000000000000000000000000000000000000",--1
								    "0000000000000000000000000000000000000000",--2
								    "0000000000000000000000000000000000000000",--3
								    "0000000000000000000000000000000000000000",--4
									 "0000000000000000000000000000000000000000",--5
									 "0000000000000000000000000000000000000000",--6
									 "0000000000000000000000000000000000000000",--7
									 "0000000000000000000000000000000000000000",--8
									 "0000000000000000000000000000000000000000",--9
								    "0000000000000000000000000000000000000000",--10         --iki nokta
								    "0000000000000000000000000000000000000000",--11
								    "0000000000000000000000000000000000000000",--12
								    "0000000000000000000000000000000000000000",--13
								    "0000000000000000000000000000000000000000",--14
								    "0000000000111111111111111111110000000000",--15
								    "0000000000111111111111111111110000000000",--16
								    "0000000000111111111111111111110000000000",--17
								    "0000000000111111111111111111110000000000",--18
								    "0000000000111111111111111111110000000000",--19
								    "0000000000111111111111111111110000000000",     --20
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000");
									 
--internal signals:: yukarıya al sonra...
signal hour_check	: integer;
	

begin

--shift the clock to left, right up and down 
	process(GPIO_0(0), GPIO_0(1), GPIO_0(2),clk_low)
	begin
		if(rising_edge(clk_low)) then
			if GPIO_0(0)='0' then
				xcoord_init_dig <= xcoord_init_dig + 1;
				xcoord_end_dig <= xcoord_end_dig + 1;
			elsif GPIO_0(1)='0' then
				xcoord_init_dig <= xcoord_init_dig - 1;
				xcoord_end_dig <= xcoord_end_dig - 1;
			elsif GPIO_0(2)='0' then
				ycoord_init_dig <= ycoord_init_dig + 1;
				ycoord_end_dig <= ycoord_end_dig + 1;
			elsif GPIO_0(3)='0' then
				ycoord_init_dig <= ycoord_init_dig - 1;
				ycoord_end_dig <= ycoord_end_dig - 1;
			end if;
		end if;
	end process;

	process(clk_40, hpos,vpos,videoOn)
	begin
		if rising_edge(clk_40) then
			if videoOn = '1' then
				if ((hpos >= xcoord_init_dig AND hpos < xcoord_end_dig) AND (vpos>=ycoord_init_dig AND vpos < ycoord_end_dig)) then
					hpos1_dig <= (hpos - xcoord_init_dig-1) mod 40;
					vpos1_dig <= (vpos - ycoord_init_dig);
					hpos2_dig <= (hpos - xcoord_init_dig);
				end if;
			end if;
		end if;
	end process;

--hour_check_p: process(cntr59_hour)
--begin
--	if cntr59_hour = 4 then
--		cntr59_hour_sig <= cntr59_hour_sig + 1;
--		if cntr59_hour_sig = 11 then
--			cntr59_hour_sig <= 0;
--		end if;
--	end if;
--end process;

cntr59_hour_sig <=  cntr59_hour; -- burayı düzenle.

draw:process(clk_40, hPos, vPos, videoOn)
	variable bmbit_dig: std_logic;
	variable bmbit_dig0: std_logic;
	variable bmbit_dig1: std_logic;
	variable bmbit_dig2: std_logic;
	variable bmbit_dig3: std_logic;
	variable bmbit_dig4: std_logic;
	variable bmbit_dig5: std_logic;
	variable bmbit_dig6: std_logic;
	variable bmbit_dig7: std_logic;
	variable bmbit_dig8: std_logic;
	
begin
	if(clk_40'event and clk_40 = '1')then
		if(videoOn = '1')then

			if ((hpos >= xcoord_init_dig and hpos < xcoord_end_dig) and (vpos >= ycoord_init_dig and vpos < ycoord_end_dig)) then
			
				if ((hpos2_dig >= 360 AND hpos2_dig < 400) AND (vpos1_dig >= 0 AND vpos1_dig < 80)) THEN
					bmbit_dig8:= BM_BOS_dig(vpos1_dig)(hpos1_dig);
					if bmbit_dig8='1' then
						VGA_R_sig <= "0000000000";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					else
						VGA_R_sig <= "0000000000";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					end if;
				
				elsif ((hpos2_dig >= 320 AND hpos2_dig < 360) AND (vpos1_dig >= 0 AND vpos1_dig < 80)) THEN
					if(cntr59 mod 10 = 0) then	
						bmbit_dig:= BM_0_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59 mod 10 = 1) then	
						bmbit_dig:= BM_1_dig(vpos1_dig)(hpos1_dig);	
					elsif(cntr59 mod 10 = 2) then	
						bmbit_dig:= BM_2_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59 mod 10 = 3) then	
						bmbit_dig:= BM_3_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59 mod 10 = 4) then	
						bmbit_dig:= BM_4_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59 mod 10 = 5) then	
						bmbit_dig:= BM_5_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59 mod 10 = 6) then	
						bmbit_dig:= BM_6_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59 mod 10 = 7) then	
						bmbit_dig:= BM_7_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59 mod 10 = 8) then	
						bmbit_dig:= BM_8_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59 mod 10 = 9) then	
						bmbit_dig:= BM_9_dig(vpos1_dig)(hpos1_dig);
					end if;
					
					if bmbit_dig = '1' then
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					else
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "1111111111";
						VGA_B_sig <= "1111111111";
					end if;
				
				elsif ((hpos2_dig >= 280 AND hpos2_dig < 320) AND (vpos1_dig >= 0 AND vpos1_dig < 80)) THEN
					
					if cntr59 < 10 then 
						bmbit_dig1:= BM_0_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59 < 20 then 
						bmbit_dig1:=BM_1_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59 < 30 then  
						bmbit_dig1:= BM_2_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59 < 40 then 
						bmbit_dig1:= BM_3_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59 < 50 then  
						bmbit_dig1:= BM_4_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59 <60 then  
						bmbit_dig1:= BM_5_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59 =60 then  
						bmbit_dig1:= BM_0_dig(vpos1_dig)(hpos1_dig);
					end if;
					
					if bmbit_dig1 = '1' then
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					else
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "1111111111";
						VGA_B_sig <= "1111111111";
					end if;
					
				elsif ((hpos2_dig >= 240 AND hpos2_dig < 280) AND (vpos1_dig >= 0 AND vpos1_dig < 80)) THEN
					bmbit_dig2:= BM_iki_nokta_dig(vpos1_dig)(hpos1_dig);
					if bmbit_dig2='1' then
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					else
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "1111111111";
						VGA_B_sig <= "1111111111";
					end if;
					
				--dakika için
				elsif ((hpos2_dig >= 200 AND hpos2_dig < 240) AND (vpos1_dig >= 0 AND vpos1_dig < 80)) THEN
					
					if(cntr59_min mod 10 = 0) then	
						bmbit_dig3:= BM_0_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_min mod 10 = 1) then	
						bmbit_dig3:= BM_1_dig(vpos1_dig)(hpos1_dig);	
					elsif(cntr59_min mod 10 = 2) then	
						bmbit_dig3:= BM_2_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_min mod 10 = 3) then	
						bmbit_dig3:= BM_3_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_min mod 10 = 4) then	
						bmbit_dig3:= BM_4_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_min mod 10 = 5) then	
						bmbit_dig3:= BM_5_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_min mod 10 = 6) then	
						bmbit_dig3:= BM_6_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_min mod 10 = 7) then	
						bmbit_dig3:= BM_7_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_min mod 10 = 8) then	
						bmbit_dig3:= BM_8_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_min mod 10 = 9) then	
						bmbit_dig3:= BM_9_dig(vpos1_dig)(hpos1_dig);
					end if;
					
					if bmbit_dig3 = '1' then
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					else
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "1111111111";
						VGA_B_sig <= "1111111111";
					end if;
					
				elsif ((hpos2_dig >= 160 AND hpos2_dig < 200) AND (vpos1_dig >= 0 AND vpos1_dig < 80)) THEN
					
					if cntr59_min < 10 then 
						bmbit_dig4:= BM_0_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_min < 20 then 
						bmbit_dig4:=BM_1_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_min < 30 then  
						bmbit_dig4:= BM_2_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_min < 40 then 
						bmbit_dig4:= BM_3_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_min < 50 then  
						bmbit_dig4:= BM_4_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_min <60 then  
						bmbit_dig4:= BM_5_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_min =60 then  
						bmbit_dig4:= BM_0_dig(vpos1_dig)(hpos1_dig);
					end if;
					
					if bmbit_dig4 = '1' then
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					else
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "1111111111";
						VGA_B_sig <= "1111111111";
					end if;
					
					
				elsif ((hpos2_dig >= 120 AND hpos2_dig < 160) AND (vpos1_dig >= 0 AND vpos1_dig < 80)) THEN
					bmbit_dig5:= BM_iki_nokta_dig(vpos1_dig)(hpos1_dig);
					if bmbit_dig5 = '1' then
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					else
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "1111111111";
						VGA_B_sig <= "1111111111";
					end if;
					
				--for hours
				elsif ((hpos2_dig >= 80 AND hpos2_dig < 120) AND (vpos1_dig >= 0 AND vpos1_dig < 80)) THEN
					
					if(cntr59_hour_sig mod 10 = 0) then	
						bmbit_dig6:= BM_0_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_hour_sig mod 10 = 1) then	
						bmbit_dig6:= BM_1_dig(vpos1_dig)(hpos1_dig);	
					elsif(cntr59_hour_sig mod 10 = 2) then	
						bmbit_dig6:= BM_2_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_hour_sig mod 10 = 3) then	
						bmbit_dig6:= BM_3_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_hour_sig mod 10 = 4) then	
						bmbit_dig6:= BM_4_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_hour_sig mod 10 = 5) then	
						bmbit_dig6:= BM_5_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_hour_sig mod 10 = 6) then	
						bmbit_dig6:= BM_6_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_hour_sig mod 10 = 7) then	
						bmbit_dig6:= BM_7_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_hour_sig mod 10 = 8) then	
						bmbit_dig6:= BM_8_dig(vpos1_dig)(hpos1_dig);
					elsif(cntr59_hour_sig mod 10 = 9) then	
						bmbit_dig6:= BM_9_dig(vpos1_dig)(hpos1_dig);
					end if;
					
					if bmbit_dig6 = '1' then
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					else
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "1111111111";
						VGA_B_sig <= "1111111111";
					end if;
					
					
				elsif ((hpos2_dig >= 40 AND hpos2_dig < 80) AND (vpos1_dig >= 0 AND vpos1_dig < 80)) THEN
					
					if cntr59_hour_sig < 10 then 
						bmbit_dig7:= BM_0_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_hour_sig < 20 then 
						bmbit_dig7:=BM_1_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_hour_sig < 30 then  
						bmbit_dig7:= BM_2_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_hour_sig < 40 then 
						bmbit_dig7:= BM_3_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_hour_sig < 50 then  
						bmbit_dig7:= BM_4_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_hour_sig <60 then  
						bmbit_dig7:= BM_5_dig(vpos1_dig)(hpos1_dig);
					elsif cntr59_hour_sig =60 then  
						bmbit_dig7:= BM_0_dig(vpos1_dig)(hpos1_dig);
					end if;
					
					if bmbit_dig7 = '1' then
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					else
						VGA_R_sig <= "1111111111";
						VGA_G_sig <= "1111111111";
						VGA_B_sig <= "1111111111";
					end if;
					
				elsif ((hpos2_dig >= 0 AND hpos2_dig < 40) AND (vpos1_dig >= 0 AND vpos1_dig < 80)) THEN
					bmbit_dig0:= BM_BOS_dig(vpos1_dig)(hpos1_dig);
					if bmbit_dig0='1' then
						VGA_R_sig <= "0000000000";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					else
						VGA_R_sig <= "0000000000";
						VGA_G_sig <= "0000000000";
						VGA_B_sig <= "0000000000";
					end if;
						
				else
					VGA_R_sig <= "1111111111";
					VGA_G_sig <= "0000000000";
					VGA_B_sig <= "1111111111";
	
				end if;
				
			else
				VGA_R_sig <= "0000000000";
			   VGA_G_sig <= "0000000000";
				VGA_B_sig <= "0000000000";
				
			end if;
			
		else
			VGA_R_sig <= "0000000000";
			VGA_G_sig <= "0000000000";
			VGA_B_sig <= "0000000000";
		end if;
	end if;
end process;

VGA_R <= VGA_R_sig;
VGA_G <= VGA_G_sig;
VGA_B <= VGA_B_sig;



end architecture;